spice


.model pch pmos(
+level=2)

.list
.end
